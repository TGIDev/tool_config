// <description>
always_comb
begin : always_comb_name
    // Combinatory
end

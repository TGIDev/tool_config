//////////////////////////////////////////////////////////////////////////////////////-
//     _____   ______    _____   _    _   _____    ______            _____    _____
//    / ____| |  ____|  / ____| | |  | | |  __ \\  |  ____|          |_   _|  / ____|
//   | (___   | |__    | |      | |  | | | |__) | | |__     ______    | |   | |
//    \\___ \\  |  __|   | |      | |  | | |  _  /  |  __|   |______|   | |   | |
//    ____) | | |____  | |____  | |__| | | | \\ \\  | |____            _| |_  | |____
//   |_____/  |______|  \\_____|  \\____/  |_|  \\_\\ |______|          |_____|  \\_____|
//
//////////////////////////////////////////////////////////////////////////////////////-
// © Copyright $CURRENT_YEAR Secure-IC S.A.S.
// This file is part of SIC-Trusted IP cores family from Secure-IC S.A.S.
// This file relies on Secure-IC S.A.S. patent portfolio.
// This file cannot be used nor duplicated without prior approval from Secure-IC S.A.S.
//////////////////////////////////////////////////////////////////////////////////////-
// Product: 
// Entity:
// File:
// Author:
// Description:

//////////////////////////////////////////////////////////////////////////////

module //Module name
#(
    // parameter Generic = x,
)(
    input logic clk,
    input logic rst_n,
);

endmodule

case ()
    val_1   :   // val = ;
    default :   // val = 
endcase
